`ifndef TYPEDEFS
`define TYPEDEFS

typedef logic [63:0] r64;
typedef logic [31:0] r32;
typedef logic [15:0] r16;
typedef logic [7:0] r8;
typedef logic [63:0] w64;
typedef logic [31:0] w32;
typedef logic [16:0] w16;
typedef logic [7:0] w8;
typedef logic [63:0] u64;
typedef logic [31:0] u32;
typedef logic [15:0] u16;
typedef logic [7:0] u8;

`endif  // TYPEDEFS