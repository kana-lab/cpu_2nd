typedef reg [31:0] r32;
typedef reg [7:0] r8;
typedef wire [31:0] w32;
typedef wire [7:0] w8;
